---bitwise 4-BIT ALU
Library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ALU4 is
PORT
 (
	 A, B		: IN STD_LOGIC_VECTOR(3 DOWNTO 0); --ONE BIT CONTROL WHICH WILL BE THE 3RD BIT OF THE SEL FOR THE ALU 
	 SEL			: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	 CIN, LESS	: IN STD_LOGIC;
	 F				: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	 COUT, OVERFLOW, SET, ZERO	: OUT STD_LOGIC
 );
END ALU4;

architecture ARCH of ALU4  is
COMPONENT ADD4
PORT
 (
	 x_in, Y_in	: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	 carry_in1 	: IN STD_LOGIC;
	 sum 			: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	 carry_out 	: OUT STD_LOGIC
 );
END COMPONENT;

COMPONENT BWOR4
--BWOR4 PORT GOES HERE
PORT
 (
	 x_IN, Y_IN 		: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	 Z_OUT		: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)	
 );
END COMPONENT;

COMPONENT BWAND4
--BWAND4 PORT GOES HERE
PORT
 (
	 x_IN , Y_IN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	 Z_OUT		: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)	
 );
END COMPONENT;

COMPONENT PINV4
--BWINV4 PORT GOES HERE
PORT
 (
	 x_IN 		: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	 y_OUT		: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SEL			: IN STD_LOGIC -- ONE BIT CONTROL WHICH WILL BE THE 3RD BIT OF THE SEL FOR THE ALU
 );
END COMPONENT;

COMPONENT MUX4X4
PORT(
	w0,w1,w2,w3 : IN STD_LOGIC_Vector(3 DOWNTO 0); -- 4 4-bit inputs
		S			: IN STD_LOGIC_Vector(1 DOWNTO 0);
		f			: OUT STD_LOGIC_Vector(3 DOWNTO 0));
END COMPONENT;

-- signals goes here
	SIGNAL ADDOUT,OROUT,ANDOUT,INVOUT,SLTOUT,MUXOUT : STD_LOGIC_Vector(3 DOWNTO 0);
	SIGNAL LESSMUX :STD_LOGIC_Vector(3 DOWNTO 0);
BEGIN
--portmap goes here

AND1: BWAND4 PORT MAP(A, B, ANDOUT);
OR1: BWOR4 PORT MAP(A, B, OROUT);
IN1: PINV4 PORT MAP(B, INVOUT, SEL(2));
ADDER1: ADD4 PORT MAP(A, INVOUT, CIN,ADDOUT,COUT); -- THIS WILL ALSO BE USED FOR SUBTRACTION
MUX1: MUX4X4 PORT MAP(ANDOUT,OROUT,ADDOUT,LESSMUX, SEL(1 DOWNTO 0),MUXOUT); --AND=00, OR=01, ADD/SUBTRACT=10, SLT = 11

--For the least significant bit Less value should be sign of A – B
PROCESS(A,B,LESS,CIN,SEL)
BEGIN

F <= MUXOUT;
OVERFLOW <= (NOT A(3) AND NOT INVOUT(3) AND ADDOUT(3)) OR (A(3) AND INVOUT(3) AND NOT ADDOUT(3));
--Overflow <= A(3) AND B(3); -- CHECKS TO SEE IF BOTH OF THE MSB ARE 1, THIS WILL CAUSE AN OVERFLOW
LESSMUX <= ("000" & LESS); --A + ~B + 1= A-B
SET <= ADDOUT(3);--(A(3) OR NOT B(3) OR '1');
ZERO <= ADDOUT(3) OR ADDOUT(2) OR ADDOUT(1) OR ADDOUT(0); -- THESE ARE ORING THE RESULTS FROM EACH ALU, AT THE END "OR" ALL ZEROS AND NEGATE



	 END PROCESS;
END ARCH;