Library IEEE;
use ieee.std_logic_1164.all;

ENTITY MUXTEST IS
PORT(
		Q0,Q1,Q2,Q3,Q4,Q5,Q6,Q7	: IN STD_LOGIC_Vector(15 DOWNTO 0);--THESE WILL BE 8 BIT INPUT FROM THE REGISTERS
		S									: IN STD_LOGIC_Vector(2 DOWNTO 0); --SELECT BIT, WE HAVE 3 BITS OF INPUT BUT ARE ONLY USING THE FIRST TWO BITS 
		FOUT_1							: OUT STD_LOGIC_Vector(15 DOWNTO 0)); --THIS IS WHAT WILL BE OUTPUT FROM THE GIANT MUX
		--BELOW HERE IS FOR THE SECOND ADDRESS TO BE READ
--		Q2_0,Q2_1,Q2_2,Q2_3,Q2_4,Q2_5,Q2_6,Q2_7	: IN STD_LOGIC_Vector(15 DOWNTO 0);--THESE WILL BE 8 BIT INPUT FROM THE REGISTERS
--		S2															: IN STD_LOGIC_Vector(2 DOWNTO 0); --SELECT BIT, WE HAVE 3 BITS OF INPUT BUT ARE ONLY USING THE FIRST TWO BITS 
--		FOUT_2													: OUT STD_LOGIC_Vector(15 DOWNTO 0)); --THIS IS WHAT WILL BE OUTPUT FROM THE GIANT MUX

END ENTITY;
ARCHITECTURE STRUCT OF MUXTEST IS 

	COMPONENT MUX4X4 IS
	PORT(
		w0,w1,w2,w3 : IN STD_LOGIC_Vector(3 DOWNTO 0); -- 4 bit input? does this mean the output will need to be a STD vector too?
			S			: IN STD_LOGIC_Vector(1 DOWNTO 0);
			f			: OUT STD_LOGIC_Vector(3 DOWNTO 0));
	
	END COMPONENT;

SIGNAL M1OUT_1,M1OUT_2,M1OUT_3,M1OUT_4 : STD_LOGIC_Vector(3 DOWNTO 0);
SIGNAL M2OUT_1,M2OUT_2,M2OUT_3,M2OUT_4 : STD_LOGIC_Vector(3 DOWNTO 0);
SIGNAL M3OUT : STD_LOGIC_Vector(15 DOWNTO 0);
-- bELOW HERE IS FOR THE SECOND REGISTER ADDRESS
--SIGNAL M2_1OUT_1,M2_1OUT_2,M2_1OUT_3,M2_1OUT_4 : STD_LOGIC_Vector(3 DOWNTO 0);
--SIGNAL M2_2OUT_1,M2_2OUT_2,M2_2OUT_3,M2_2OUT_4 : STD_LOGIC_Vector(3 DOWNTO 0);
--SIGNAL M2_3OUT : STD_LOGIC_Vector(15 DOWNTO 0);
BEGIN 


QOUT0 : MUX4X4 PORT MAP(Q0(3 DOWNTO 0),Q1(3 DOWNTO 0),Q2(3 DOWNTO 0),Q3(3 DOWNTO 0),S(1 DOWNTO 0),M1OUT_1); --M1OUT [3..0]
QOUT1 : MUX4X4 PORT MAP(Q0(7 DOWNTO 4),Q1(7 DOWNTO 4),Q2(7 DOWNTO 4),Q3(7 DOWNTO 4),S(1 DOWNTO 0),M1OUT_2);--M1OUT [7..4]
QOUT2 : MUX4X4 PORT MAP(Q0(11 DOWNTO 8),Q1(11 DOWNTO 8),Q2(11 DOWNTO 8),Q3(11 DOWNTO 8),S(1 DOWNTO 0),M1OUT_3);--M1OUT [11..8]
QOUT3 : MUX4X4 PORT MAP(Q0(15 DOWNTO 12),Q1(15 DOWNTO 12),Q2(15 DOWNTO 12),Q3(15 DOWNTO 12),S(1 DOWNTO 0),M1OUT_4);--M1OUT [15..12]


QOUT4 : MUX4X4 PORT MAP(Q4(3 DOWNTO 0),Q5(3 DOWNTO 0),Q6(3 DOWNTO 0),Q7(3 DOWNTO 0),S(1 DOWNTO 0),M2OUT_1);--M2OUT [3..0]
QOUT5 : MUX4X4 PORT MAP(Q4(7 DOWNTO 4),Q5(7 DOWNTO 4),Q6(7 DOWNTO 4),Q7(7 DOWNTO 4),S(1 DOWNTO 0),M2OUT_2); --M2OUT [7..4]
QOUT6 : MUX4X4 PORT MAP(Q4(11 DOWNTO 8),Q5(11 DOWNTO 8),Q6(11 DOWNTO 8),Q7(11 DOWNTO 8),S(1 DOWNTO 0),M2OUT_3); --M2OUT [11..8]
QOUT7 : MUX4X4 PORT MAP(Q4(15 DOWNTO 12),Q5(15 DOWNTO 12),Q6(15 DOWNTO 12),Q7(15 DOWNTO 12),S(1 DOWNTO 0),M2OUT_4); --M2OUT [15..12]


QOUT_3_0 : MUX4X4 PORT MAP(M1OUT_1,M1OUT_1,M2OUT_1,M2OUT_1,S(2 DOWNTO 1),M3OUT(3 DOWNTO 0));
QOUT_7_4 : MUX4X4 PORT MAP(M1OUT_2,M1OUT_2,M2OUT_2,M2OUT_2,S(2 DOWNTO 1),M3OUT(7 DOWNTO 4));
QOUT_11_8 : MUX4X4 PORT MAP(M1OUT_3,M1OUT_3,M2OUT_3,M2OUT_3,S(2 DOWNTO 1),M3OUT(11 DOWNTO 8));
QOUT_15_12 : MUX4X4 PORT MAP(M1OUT_4,M1OUT_4,M2OUT_4,M2OUT_4,S(2 DOWNTO 1),M3OUT(15 DOWNTO 12));
FOUT_1<=M3OUT;

-- BELOW HERE IS FOR THE SECOND REGISTER ADDRESS TO BE READ

--Q2_OUT0 : MUX4X4 PORT MAP(Q2_0(3 DOWNTO 0),Q2_1(3 DOWNTO 0),Q2_2(3 DOWNTO 0),Q2_3(3 DOWNTO 0),S2(1 DOWNTO 0),M2_1OUT_1); --M2_1OUT [3..0]
--Q2_OUT1 : MUX4X4 PORT MAP(Q2_0(7 DOWNTO 4),Q2_1(7 DOWNTO 4),Q2_2(7 DOWNTO 4),Q2_3(7 DOWNTO 4),S2(1 DOWNTO 0),M2_1OUT_2);--M2_1OUT [7..4]
--Q2_OUT2 : MUX4X4 PORT MAP(Q2_0(11 DOWNTO 8),Q2_1(11 DOWNTO 8),Q2_2(11 DOWNTO 8),Q2_3(11 DOWNTO 8),S2(1 DOWNTO 0),M2_1OUT_3);--M2_1OUT [11..8]
--Q2_OUT3 : MUX4X4 PORT MAP(Q2_0(15 DOWNTO 12),Q2_1(15 DOWNTO 12),Q2_2(15 DOWNTO 12),Q2_3(15 DOWNTO 12),S2(1 DOWNTO 0),M2_1OUT_4);--M2_1OUT [15..12]
--
--
--Q2_OUT4 : MUX4X4 PORT MAP(Q2_4(3 DOWNTO 0),Q2_5(3 DOWNTO 0),Q2_6(3 DOWNTO 0),Q2_7(3 DOWNTO 0),S2(1 DOWNTO 0),M2_2OUT_1);--M2_2OUT [3..0]
--Q2_OUT5 : MUX4X4 PORT MAP(Q2_4(7 DOWNTO 4),Q2_5(7 DOWNTO 4),Q2_6(7 DOWNTO 4),Q2_7(7 DOWNTO 4),S2(1 DOWNTO 0),M2_2OUT_2); --M2_2OUT [7..4]
--Q2_OUT6 : MUX4X4 PORT MAP(Q2_4(11 DOWNTO 8),Q2_5(11 DOWNTO 8),Q2_6(11 DOWNTO 8),Q2_7(11 DOWNTO 8),S2(1 DOWNTO 0),M2_2OUT_3); --M2_2OUT [11..8]
--Q2_OUT7 : MUX4X4 PORT MAP(Q2_4(15 DOWNTO 12),Q2_5(15 DOWNTO 12),Q2_6(15 DOWNTO 12),Q2_7(15 DOWNTO 12),S2(1 DOWNTO 0),M2_2OUT_4); --M2_2OUT [15..12]
--
--
--Q2OUT_3_0 : MUX4X4 PORT MAP(M2_1OUT_1,M2_1OUT_1,M2_2OUT_1,M2_2OUT_1,S(2 DOWNTO 1),M2_3OUT(3 DOWNTO 0));
--Q2OUT_7_4 : MUX4X4 PORT MAP(M2_1OUT_2,M2_1OUT_2,M2_2OUT_2,M2_2OUT_2,S(2 DOWNTO 1),M2_3OUT(7 DOWNTO 4));
--Q2OUT_11_8 : MUX4X4 PORT MAP(M2_1OUT_3,M2_1OUT_3,M2_2OUT_3,M2_2OUT_3,S(2 DOWNTO 1),M2_3OUT(11 DOWNTO 8));
--Q2OUT_15_12 : MUX4X4 PORT MAP(M2_1OUT_4,M2_1OUT_4,M2_2OUT_4,M2_2OUT_4,S(2 DOWNTO 1),M2_3OUT(15 DOWNTO 12));
--FOUT_2<=M2_3OUT;


END STRUCT;