--ADD16
--Design a 16-bit adding machine, ADD16 (using ADD4)
Library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ADD16 is
PORT
 (
	 x_in, Y_in	: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	 carry_in1 	: IN STD_LOGIC;
	 sum 			: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	 carry_out 	: OUT STD_LOGIC
 );

END ADD16;

architecture STRUCT OF ADD16 IS 
--COMPONENTS HERE 
COMPONENT ADD4 IS 
PORT
 (
	 x_in, Y_in	: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	 carry_in1 	: IN STD_LOGIC;
	 sum 			: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	 carry_out 	: OUT STD_LOGIC
 );
END COMPONENT;
--SIGNALS HERE 
SIGNAL CARRY_OUT_VECTOR : STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN

--PORTMAPS HERE	
ADD0: ADD4 PORT MAP(x_in(3 DOWNTO 0),Y_in(3 DOWNTO 0),CARRY_IN1,SUM(3 DOWNTO 0),CARRY_OUT_VECTOR(0));
ADD1: ADD4 PORT MAP(x_in(7 DOWNTO 4),Y_in(7 DOWNTO 4),CARRY_OUT_VECTOR(0),SUM(7 DOWNTO 4),CARRY_OUT_VECTOR(1));
ADD2: ADD4 PORT MAP(x_in(11 DOWNTO 8),Y_in(11 DOWNTO 8),CARRY_OUT_VECTOR(1),SUM(11 DOWNTO 8),CARRY_OUT_VECTOR(2));
ADD3: ADD4 PORT MAP(x_in(15 DOWNTO 12),Y_in(15 DOWNTO 12),CARRY_OUT_VECTOR(2),SUM(15 DOWNTO 12),CARRY_OUT_VECTOR(3));

CARRY_OUT <= CARRY_OUT_VECTOR(3);
--PROCESS HERE

END STRUCT;